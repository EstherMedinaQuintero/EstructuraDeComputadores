/// Podemos definir constantes en verilog
/// Y al instanciar podemos poner un valor distinto

module mux2 #(parameter WIDTH = 8) (output wire [WIDTH-1:0], blabla)
endmodule

/// #retardo

/// Máquina de estados finitos
  /// ¿Qué quiero?
  /// ¿Qué estados?
    /// Dónde transito
    /// Con qué salida
/// Contador de unos (EJEMPLO)
  /// Siempre miramos el menos significativo